module riscv_cpu_core(

);

endmodule
