module riscv_cpu_fetch_unit(

);

endmodule

