module riscv_cpu_exec_unit(

);

endmodule
