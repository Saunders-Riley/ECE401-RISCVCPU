module riscv_cpu_integration(

);

endmodule
