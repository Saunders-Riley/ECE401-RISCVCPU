module riscv_cpu_commit_unit(

);

endmodule
